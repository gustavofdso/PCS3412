-- PCS3412 - Organizacao e Arquitetura de Computadores I
-- Project: T-FIVE-MC
-- File: FD.vhd
-- Author: Gustavo Freitas de Sá Oliveira
--
-- Description:
--     Contém o fluxo de dados, com todos os seus componentes ligados

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.constants.all;
use work.types.all;
